module gal2 ( 
	clk,
	clr,
	lb,
	eb,
	ec,
	disp
	) ;

input  clk;
input  clr;
input  lb;
input  eb;
input  ec;
inout [6:0] disp;
