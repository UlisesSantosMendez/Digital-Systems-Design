module contador ( 
	clk,
	en,
	clr,
	q
	) ;

input  clk;
input  en;
inout  clr;
inout [9:0] q;
