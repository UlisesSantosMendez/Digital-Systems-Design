module contador ( 
	clk,
	clr,
	sen,
	uni,
	dec
	) ;

input  clk;
input  clr;
input [1:0] sen;
inout [3:0] uni;
inout [2:0] dec;
