module mensaje ( 
	clr,
	clk,
	display,
	cat
	) ;

input  clr;
input  clk;
inout [6:0] display;
inout [2:0] cat;
