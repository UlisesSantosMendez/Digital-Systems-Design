module gal1 ( 
	clk,
	clr,
	ini,
	z,
	a0,
	ec,
	eb,
	lb,
	la,
	ea
	) ;

input  clk;
input  clr;
input  ini;
input  z;
input  a0;
inout  ec;
inout  eb;
inout  lb;
inout  la;
inout  ea;
