module mealy ( 
	clk,
	clr,
	e,
	dis
	) ;

input  clk;
input  clr;
inout  e;
inout [6:0] dis;
