module marq ( 
	clk,
	clr,
	e,
	display
	) ;

input  clk;
input  clr;
input [2:0] e;
inout [9:0] display;
