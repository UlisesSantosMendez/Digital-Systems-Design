module mealy ( 
	clk,
	clr,
	e,
	s,
	dis
	) ;

input  clk;
input  clr;
input  e;
inout  s;
inout [6:0] dis;
