module gal1 ( 
	clk,
	clr,
	ini,
	d,
	ec,
	eb,
	lb,
	a
	) ;

input  clk;
input  clr;
input  ini;
input [5:0] d;
inout  ec;
inout  eb;
inout  lb;
inout [5:0] a;
