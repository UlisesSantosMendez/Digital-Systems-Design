module counter ( 
	clk,
	clr,
	en,
	q
	) ;

input  clk;
input  clr;
input  en;
inout [2:0] q;
