module boleta ( 
	clk,
	clr,
	en,
	display
	) ;

input  clk;
input  clr;
input  en;
inout [6:0] display;
