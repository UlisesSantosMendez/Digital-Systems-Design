module contador ( 
	clk,
	clr,
	en,
	q
	) ;

input  clk;
input  clr;
input  en;
inout [9:0] q;
